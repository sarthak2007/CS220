`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:50:50 01/21/2019 
// Design Name: 
// Module Name:    two-bit-adder 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module two_bit_adder(x,y,z,carry
    );
input [1:0] x;
input [1:0] y;
output [1:0] z;
wire [1:0] z;
output carry;
wire carry ;
wire carry0;

endmodule
